module testbench;

    parameter WIDTH=32;
    parameter PERIOD=20;

    logic clk, rst_n;
    // tb - master wire
    wire [WIDTH-1 : 0]  tb_master_data;
    wire                tb_master_valid;
    wire                master_tb_ready;
    // master - slave wire
    wire [WIDTH-1 : 0]  master_slave_data;
    wire                master_slave_valid;
    wire                slave_master_ready;
    // slave - tb wire
    wire [WIDTH-1 : 0]  slave_tb_data;
    wire                slave_tb_valid;
    wire                tb_slave_ready;

    node(.WIDTH(WIDTH)) master(
                            //input 
                            .clk(clk), 
                            .rst_n(rst_n),
                            .data_in(tb_master_data),
                            .valid_up_in(tb_master_valid), 
                            .ready_down_in(slave_master_ready),
                            //output
                            .data_out(master_slave_data),
                            .valid_down_out(master_slave_valid),
                            .ready_up_out(master_tb_ready)
                        );

    node(.WIDTH(WIDTH)) slave(
                            //input 
                            .clk(clk), 
                            .rst_n(rst_n),
                            .data_in(master_slave_data),
                            .valid_up_in(master_slave_valid), 
                            .ready_down_in(tb_slave_ready),
                            //output
                            .data_out(slave_tb_data),
                            .valid_down_out(slave_tb_valid),
                            .ready_up_out(slave_master_ready)
                        );

    always #(PERIOD/2) clk = ~clk;

    initial begin
        #1
        $dumpfile("wave.vcd");
		$dumpvars;
        clk             = 1'b1;
        rst_n           = 1'b0;
        tb_slave_ready  = 1'b0;
        tb_master_valid = 1'b0;

        repeat (10) @(posedge clk);
        rst_n           = 1'b1;
        tb_slave_ready  = 1'b1;
        tb_master_valid = 1'b1;

        //TODO: task for vld-invalid-valid pattern

        //TODO: task for sequential pattern

        
    end
    
endmodule